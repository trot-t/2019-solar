boost converter
.MODEL swmod SW(Roff=1000000 Ron=1 VT=.98 VH=.001)
V1 1 0 85
L1 1 2 0.102
lk 2 2a 1p    ;current transformer for mesurement 
lr 3 3a 1p    ;current transformer
D1 2 3 D
C1 3 0 0.75uF
R1 3a 0 1157.76
SW 2a 0 ns1 0 swmod 
VS1 ns1 0 PWL(0 0 .1m 0 .1m 1 .2m 1 .2m 0) R=0
.control
tran .001m 14m 
plot V(1), V(3)
plot L1#branch,lr#branch
* gnuplot boost_result V(1),V(3)
.endc
.end
